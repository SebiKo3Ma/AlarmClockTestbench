class scoreboard_queues;
    config_transaction cfg[$];
    alarm_transaction  al[$];
endclass