package config_pkg;
    int verbosity = 0;  // Default verbosity level
    string test_name;
endpackage
