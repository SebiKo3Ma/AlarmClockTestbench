typedef enum logic[1:0]{
  CR,
  OP,
  AL,
  IL} trans_types;
