package config_pkg;
    int verbosity = 0;  // Default verbosity level
endpackage
